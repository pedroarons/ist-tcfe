ngspice T2-1 
 
.options savecurrents 
 
Vs n1 GND 5.178860 
V0 GND n9 0 
R1 n2 n1 1.023629k 
R2 n3 n2 2.086404k 
R3 n2 n5 3.099961k 
R4 n5 GND 4.081833k 
R5 n6 n5 3.041696k 
R6 n7 n9 2.041567k 
R7 n8 n7 1.041568k 
H1 n5 n8 V0 8.168406k 
G1 n6 n3 n2 n5 7.295719m 
C1 n6 n8 1.049083u 
 
.control 
 
op 
echo "t2-1_TAB" 
print all 
echo "t2-1_END" 
 
quit 
.endc 
 
.end